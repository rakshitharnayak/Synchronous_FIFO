//////////////////////////////////////////////////////////////////////////
`define DATA_W 128           // Data width
`define DEPTH 1024        // Depth of FIFO
`define UPP_TH 4           // Upper threshold to generate Almost-full
`define LOW_TH 2           //  Lower threshold to generate Almost-empty
// `define ADDRESS 10
//////////////////////////////////////////////////////////////////////////
